LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

LIBRARY LPM;
USE LPM.LPM_COMPONENTS.ALL;

ENTITY ADC_INTERFACE IS
PORT(
	ADC_WCLK    : IN  STD_LOGIC;
	ADC_BCLK    : IN  STD_LOGIC;
	ADC_DAT     : IN  STD_LOGIC;
	CPU_CLK     : IN  STD_LOGIC;
	SOUND_DATA  : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	NEW_SAMPLE  : OUT STD_LOGIC
	);
END ADC_INTERFACE;

ARCHITECTURE a OF ADC_INTERFACE IS

	-- Declare signals
	signal shifted_data          : std_logic_vector(15 downto 0); -- Shift register output
	signal buffer_data           : std_logic_vector(15 downto 0); -- Output buffer
	signal write_req, read_req   : std_logic;  -- FIFO control signals
	signal rdempty, rdempty_delay : std_logic; -- New data indication
	signal bit_count             : integer range 0 to 18;   -- Counter for number of bits shifted in

BEGIN

	-- Shift register to parallelize the data from the ADC
	serialize : lpm_shiftreg
	GENERIC MAP (
		lpm_direction => "LEFT",
		lpm_type => "LPM_SHIFTREG",
		lpm_width => 16
	)
	PORT MAP (
		clock => ADC_BCLK, -- Latch data on falling edges
		q => shifted_data,      -- Output of shift register
		shiftin => ADC_DAT      -- Input to shift register
	);

	
	-- A dual-clock FIFO to ensure timing safety across clock domains
	ADC_FIFO_inst : work.ADC_FIFO PORT MAP (
		data => shifted_data,   -- Data input to the FIFO
		rdclk => CPU_CLK,       -- Read clock (synchronous to CPU_CLK)
		rdreq => read_req,      -- Read request (generated by FIFO control logic)
		wrclk => ADC_BCLK,      -- Write clock (synchronous to ADC_BCLK)
		wrreq => write_req,     -- Write request (generated by FIFO control logic)
		q => SOUND_DATA,       -- Data output from the FIFO
		rdempty => rdempty  -- Empty flag (indicates whether FIFO is empty)
	);

	
	-- Whenever new data is available, pull it out of the FIFO.
	read_req <= not rdempty;
	-- Indicate new data after data updates
	read_indication : process(CPU_CLK)
	begin
		-- Using the falling edge keeps changes away from sample times
		-- in your peripheral.  This isn't a good practice because it can
		-- cut your effective max frequency in half, but this isn't a
		-- bleeding-edge system and this is much easier than trying to
		-- design around timing constraints.
		if falling_edge(CPU_CLK) then
			-- Indicate data new after pulled from FIFO.
			rdempty_delay <= not rdempty;
			NEW_SAMPLE <= rdempty_delay;
		end if;
	end process;
	


	-- Track the number of bits coming it, and latch into FIFO when needed.
	write_control : process(ADC_BCLK)
	begin
		if rising_edge(ADC_BCLK) then
			-- Start counting when word clock is high
			if ADC_WCLK = '1' then
				bit_count <= 16;
			elsif bit_count /= 0 then
				bit_count <= bit_count - 1;
			end if;
			if bit_count = 1 then
			-- Write data to FIFO after 16 bits have been shifted in
				write_req <= '1';
			else
				write_req <= '0';
			end if;
		end if;
	end process;    
END a;
